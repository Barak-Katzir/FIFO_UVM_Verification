
`ifndef DATA_WIDTH
`define DATA_WIDTH 8
`endif

// default FIFO depth is 2^4=16 words
`ifndef ADDR_WIDTH
`define ADDR_WIDTH 4
`endif


// 2**`ADDR_WIDTH - 1